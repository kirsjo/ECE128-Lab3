`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 09/19/2023 02:56:30 PM
// Design Name: 
// Module Name: fourBitAdder_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module fourBitAdder_tb();
    reg [3:0] A, B;
    reg CI;
    wire [3:0] SUM;
    wire CO;
    
    
    fourBit uut(.A(A), .B(B), .CI(CI), .SUM(SUM), .CO(CO));
    
    
    initial begin
        A = 4'b0000; B=4'b0000; CI=0;
        #10
        A = 4'b0001; B=4'b0000;CI=0;
        #10
        A = 4'b0010; B=4'b0000;CI=0;
        #10
        A = 4'b0011; B=4'b0000;CI=0;
        #10
        A = 4'b0100; B=4'b0000;CI=0;
        #10
        A = 4'b0101; B=4'b0000;CI=0;
        #10
        A = 4'b0110; B=4'b0000;CI=0;
        #10
        A = 4'b0111; B=4'b0000;CI=0;
        #10
        A = 4'b1000; B=4'b0000;CI=0;
        #10
        A = 4'b1001; B=4'b0000;CI=0;
        #10
        A = 4'b1010; B=4'b0000;CI=0;
        #10
        A = 4'b1011; B=4'b0000;CI=0;
        #10
        A = 4'b1100; B=4'b0000; CI=0;
        #10
        A = 4'b1101; B=4'b0000;CI=0;
        #10
        A = 4'b1110; B=4'b0000;CI=0;
        #10
        A = 4'b1111; B=4'b0000;CI=0;
        #10
        A = 4'b0001; B=4'b0001;CI=0;
        #10
        A = 4'b0010; B=4'b0001;CI=0;
        #10
        A = 4'b0011; B=4'b0001;CI=0;
        #10
        A = 4'b0100; B=4'b0001;CI=0;
        #10
        A = 4'b0101; B=4'b0001;CI=0;
        #10
        A = 4'b0110; B=4'b0001;CI=0;
        #10
        A = 4'b0111; B=4'b0001;CI=0;
        #10
        A = 4'b1000; B=4'b0001;CI=0;
        #10
        A = 4'b1001; B=4'b0001;CI=0;
        #10
        A = 4'b1010; B=4'b0001;CI=0;
        #10
        A = 4'b1011; B=4'b0001;CI=0;
        #10
        A = 4'b1100; B=4'b0001;CI=0;
        #10
        A = 4'b1101; B=4'b0001;CI=0;
        #10
        A = 4'b1110; B=4'b0001;CI=0;
        #10
        A = 4'b1111; B=4'b0001;CI=0;
        #10
        A = 4'b0010; B=4'b0010;CI=0;
        #10
        A = 4'b0011; B=4'b0010;CI=0;
        #10
        A = 4'b0100; B=4'b0010;CI=0;
        #10
        A = 4'b0101; B=4'b0010;CI=0;
        #10
        A = 4'b0110; B=4'b0010;CI=0;
        #10
        A = 4'b0111; B=4'b0010;CI=0;
        #10
        A = 4'b1000; B=4'b0010;CI=0;
        #10
        A = 4'b1001; B=4'b0010;CI=0;
        #10
        A = 4'b1010; B=4'b0010;CI=0;
        #10
        A = 4'b1011; B=4'b0010;CI=0;
        #10
        A = 4'b1100; B=4'b0010;CI=0;
        #10
        A = 4'b1101; B=4'b0010;CI=0;
        #10
        A = 4'b1110; B=4'b0010;CI=0;
        #10
        A = 4'b1111; B=4'b0010;CI=0;
        #10
        A = 4'b0011; B=4'b0011;CI=0;
        #10
        A = 4'b0100; B=4'b0011;CI=0;
        #10
        A = 4'b0101; B=4'b0011;CI=0;
        #10
        A = 4'b0110; B=4'b0011;CI=0;
        #10
        A = 4'b0111; B=4'b0011;CI=0;
        #10
        A = 4'b1000; B=4'b0011;CI=0;
        #10
        A = 4'b1001; B=4'b0011;CI=0;
        #10
        A = 4'b1010; B=4'b0011;CI=0;
        #10
        A = 4'b1011; B=4'b0011;CI=0;
        #10
        A = 4'b1100; B=4'b0011;CI=0;
        #10
        A = 4'b1101; B=4'b0011;CI=0;
        #10
        A = 4'b1110; B=4'b0011;CI=0;
        #10
        A = 4'b1111; B=4'b0011;CI=0;
        #10
        A = 4'b0100; B=4'b0100;CI=0;
        #10
        A = 4'b0101; B=4'b0100;CI=0;
        #10
        A = 4'b0110; B=4'b0100;CI=0;
        #10
        A = 4'b0111; B=4'b0100;CI=0;
        #10
        A = 4'b1000; B=4'b0100;CI=0;
        #10
        A = 4'b1001; B=4'b0100;CI=0;
        #10
        A = 4'b1010; B=4'b0100;CI=0;
        #10
        A = 4'b1011; B=4'b0100;CI=0;
        #10
        A = 4'b1100; B=4'b0100;CI=0;
        #10
        A = 4'b1101; B=4'b0100;CI=0;
        #10
        A = 4'b1110; B=4'b0100;CI=0;
        #10
        A = 4'b1111; B=4'b0100;CI=0;
        #10
        A = 4'b0101; B=4'b0101;CI=0;
        #10
        A = 4'b0110; B=4'b0101;CI=0;
        #10
        A = 4'b0111; B=4'b0101;CI=0;
        #10
        A = 4'b1000; B=4'b0101;CI=0;
        #10
        A = 4'b1001; B=4'b0101;CI=0;
        #10
        A = 4'b1010; B=4'b0101;CI=0;
        #10
        A = 4'b1011; B=4'b0101;CI=0;
        #10
        A = 4'b1100; B=4'b0101;CI=0;
        #10
        A = 4'b1101; B=4'b0101;CI=0;
        #10
        A = 4'b1110; B=4'b0101;CI=0;
        #10
        A = 4'b1111; B=4'b0101;CI=0;
        #10
        A = 4'b0110; B=4'b0110;CI=0;
        #10
        A = 4'b0111; B=4'b1110;CI=0;
    end

endmodule
